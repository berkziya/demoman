module rom (
    input clk,
    input rst,
    input [9:0] addr,
    output reg [15:0] data
);

endmodule

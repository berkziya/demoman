// Transformations
//    a
//  f   b
//    g
//  e   c
//    d
//                  gfedcba
parameter _0 = 7'b1000000; // 0
parameter _1 = 7'b1111001; // 1
parameter _2 = 7'b0100100; // 2
parameter _3 = 7'b0110000; // 3
parameter _4 = 7'b0011001; // 4
parameter _5 = 7'b0010010; // 5
parameter _6 = 7'b0000010; // 6
parameter _7 = 7'b1111000; // 7
parameter _8 = 7'b0000000; // 8
parameter _9 = 7'b0010000; // 9

parameter _A = 7'b0001000; // A
parameter _B = 7'b0000011; // b
parameter _C = 7'b1000110; // C
parameter _D = 7'b0100001; // d
parameter _E = 7'b0000110; // E
parameter _F = 7'b0001110; // F
parameter _G = 7'b1000010; // G
parameter _H = 7'b0001001; // H
parameter _I = 7'b1111001; // I
parameter _J = 7'b1110001; // J
parameter _K = 7'b0001010; // (Custom K: H with a kicked leg)
parameter _L = 7'b1000111; // L
parameter _M = 7'b0101100; // (Custom M: like A with middle top, no center bar)
parameter _N = 7'b0101011; // n
parameter _O = 7'b1000000; // 0
parameter _P = 7'b0001100; // P
parameter _Q = 7'b0011000; // q
parameter _R = 7'b0101111; // r
parameter _S = 7'b0010010; // S
parameter _T = 7'b0000111; // t
parameter _U = 7'b1000001; // U
parameter _V = 7'b1100011; // (Lowercase u/v shape)
parameter _W = 7'b1000001; // (Using U for W)
parameter _X = 7'b0001001; // (Using H for X)
parameter _Y = 7'b0010001; // Y
parameter _Z = 7'b0110100; // Z

parameter _SPACE      = 7'b1111111; // ' '
parameter _DASH       = 7'b0111111; // '-'
parameter _UNDERSCORE = 7'b1110111; // '_'
parameter _LOWSQUARE  = 7'b0011100; // 'o'
parameter _HIGHSQUARE = 7'b0100011; // 'o' but flying

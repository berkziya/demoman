module hitbox ();
endmodule
